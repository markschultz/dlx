`include "./dlx.defines"

module top (clk, MRST, in, out, state, DAddr, DRead, DWrite, DOut, IRead, framebit, clkout, i);
   input clk;
	input MRST;
	input [5:0] in;
	output [15:0] out;
	output [4:0] state;
	output [3:0] i;
	
	output [`WordSize]	DAddr;          // Address for Data Cache read/write
	output					DRead;          // Data Cache read enable
	output					DWrite;         // Data Cache write enable
	output [`WordSize]	DOut;           // Data Input to Data Cache (write)
	//input  [`WordSize]	DIn;            // Data Output from Data Cache (read)
	//output [`WordSize]	IAddr;          // Instruction Cache read address
	output					IRead;          // Instruction Cache read enable
	//input  [`WordSize]	IIn;            // Instruction from Instruction Cache
	output framebit;
	output clkout;
	//output clkout1;
	
//	reg tren;
	reg [`WordSize]	IIn;
   reg [31:0] 	memory[63:0];
   wire [`WordSize] 	IAddr;
	wire [`WordSize] DIn;
	//synthesis attribute keep of i is "true";
	reg [3:0] i;
	
	assign out = IIn[15:0];
	assign DIn = {32{1'b1}};
	assign framebit = ~|(i);
	assign clkout = clk;      //&(~MRST);
	//assign clkout1 = clk;
	
	always @(negedge clk or posedge MRST) 
   begin 
		if (MRST)
		begin
			IIn <= {`SPECIAL, 5'b0, 5'b0, 5'b0, 5'b0, `NOP};
//			tren <= 1'b0;
		end
		else
		begin
			if (in[4:1] == 4'b0001) 
			begin
				IIn <= memory[i]; //IIn <= memory[((IAddr/4)%64)];
//				tren <= (i[3:2]==2'b00)?1'b1:1'b0;
			end
			else if (in[4:1] == 4'b0010)
			begin
				IIn <= memory[i+16]; //IIn <= memory[((IAddr/4)%64)];
//				tren <= (i[3:2]==2'b00)?1'b1:1'b0;
			end
			else if (in[4:1] == 4'b0100)
			begin
				IIn <= memory[i+32]; //IIn <= memory[((IAddr/4)%64)];
//				tren <= (i[3:2]==2'b00)?1'b1:1'b0;
			end
			else if (in[4:1] == 4'b1000)
			begin
				IIn <= memory[i+48]; //IIn <= memory[((IAddr/4)%64)];
//				tren <= (i[3:2]==2'b00)?1'b1:1'b0;
			end
			else
			begin
				IIn <= {`SPECIAL, 5'b0, 5'b0, 5'b0, 5'b0, `NOP};	//   NOP			
//				tren <= (i[3:2]==2'b00)?1'b1:1'b0;
			end
		end
   end
	
//	assign troin = in[0];
	assign state = in[4:0];
	assign troout = 1'b0;
//	trojan tr (.test(troin), .en(tren), .ck(clk), .troout(troout));
	
	always @(posedge clk or posedge MRST)
	begin
		if (MRST) 
			i <= 4'b0;
		else
			i <= i + 1'b1;
	end
	
	always @(posedge clk or posedge MRST)
	begin
//		memory[00] <= 32'b00000000000000000000000000100010;
//		memory[01] <= 32'b00000000000000000000100000100010;
//		memory[02] <= 32'b00000000000000000001000000100010;
//		memory[03] <= 32'b00000000000000000001100000100010;
//		memory[04] <= 32'b00000000000000000010000000100010;
//		memory[05] <= 32'b00000000000000000010100000100010;
//		memory[06] <= 32'b00000000000000000011000000100010;
//		memory[07] <= 32'b00000000000000000011100000100010;
//		memory[08] <= 32'b00000000000000000100000000100010;
//		memory[09] <= 32'b00000000000000000100100000100010;
//		memory[10] <= 32'b00000000000000000101000000100010;
//		memory[11] <= 32'b00000000000000000101100000100010;
//		memory[12] <= 32'b00000000000000000110000000100010;
//		memory[13] <= 32'b00000000000000000110100000100010;
//		memory[14] <= 32'b00000000000000000111000000100010;
//		memory[15] <= 32'b00000000000000000111100000100010;
//		memory[16] <= 32'b00000000000000001000000000100010;
//		memory[17] <= 32'b00000000000000001000100000100010;
//		memory[18] <= 32'b00000000000000001001000000100010;
//		memory[19] <= 32'b00000000000000001001100000100010;
//		memory[20] <= 32'b00000000000000001010000000100010;
//		memory[21] <= 32'b00000000000000001010100000100010;
//		memory[22] <= 32'b00000000000000001011000000100010;
//		memory[23] <= 32'b00000000000000001011100000100010;
//		memory[24] <= 32'b00000000000000001100000000100010;
//		memory[25] <= 32'b00000000000000001100100000100010;
//		memory[26] <= 32'b00000000000000001101000000100010;
//		memory[27] <= 32'b00000000000000001101100000100010;
//		memory[28] <= 32'b00000000000000001110000000100010;
//		memory[29] <= 32'b00000000000000001110100000100010;
//		memory[30] <= 32'b00000000000000001111000000100010;
//		memory[31] <= 32'b00000000000000001111100000100010;
//		memory[32] <= 32'b00100000001000010000000000000001;
//		memory[33] <= 32'b00000000001000010001000000100000;
//		memory[34] <= 32'b00000000010000100001100000100001;
//		memory[35] <= 32'b00001000000000000000000000001000;
//		memory[36] <= 32'b00000000000000000000000000000000;
//		memory[37] <= 32'b00100000001000010000000000000011;
//		memory[38] <= 32'b00000000010000010101000000101101;
//		memory[39] <= 32'b00010101010000000000000000001000;
//		memory[40] <= 32'b00000000000000000000000000000000;
//		memory[41] <= 32'b00001100000000000000000000001100;
//		memory[42] <= 32'b00000000000000000000000000000000;
//		memory[43] <= 32'b01001000100000000000000000000000;
//		memory[44] <= 32'b00000000000000000000000000000000;
//		memory[45] <= 32'b00010000010000000000000000100000;
//		memory[46] <= 32'b00000000000000000000000000000000;
//		memory[47] <= 32'b00000000010000100001000000100010;
//		memory[48] <= 32'b00100000101001010000000000110100;
//		memory[49] <= 32'b00000000000000000000000000000000;
//		memory[50] <= 32'b00000000000000000000000000000000;
//		memory[51] <= 32'b00000000000000000000000000000000;
//		memory[52] <= 32'b01001100101000000000000000000000;
//		memory[53] <= 32'b00000000000000000000000000000000;
//		memory[54] <= 32'b00000000000000000000000000000000;
//		memory[55] <= 32'b00000000000000000000000000000000;
//		memory[56] <= 32'b00000000000000000000000000000000;
//		memory[57] <= 32'b00000000000000000000000000000000;
//		memory[58] <= 32'b00000000000000000000000000000000;
//		memory[59] <= 32'b00000000000000000000000000000000;
//		memory[60] <= 32'b00000000000000000000000000000000;
//		memory[61] <= 32'b00000000000000000000000000000000;
//		memory[62] <= 32'b00000000000000000000000000000000;
//		memory[63] <= 32'b00000000000000000000000000000000;
//
//
//
//memory[00]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[01]	<=	32'b000000_00001_00001_00010_00000_100010	;
//memory[02]	<=	32'b000000_00001_00001_00011_00000_100010	;
//memory[03]	<=	32'b001111_00001_00001_10011_01100_110111	;
//memory[04]	<=	32'b001111_00010_00010_01010_11100_101001	;
//memory[05]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[06]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[07]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[08]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[09]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[10]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[11]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[12]	<=	32'b000000_00001_00010_00011_00000_100100	;
//memory[13]	<=	32'b000000_00001_00010_00011_00000_100100	;
//memory[14]	<=	32'b000000_00001_00010_00011_00000_100100	;
//memory[15]	<=	32'b000000_00001_00010_00011_00000_100100	;
//memory[16]	<=	32'b000000_00001_00010_00011_00000_100100	;
//memory[17]	<=	32'b000000_00001_00010_00011_00000_100100	;
//memory[18]	<=	32'b000000_00001_00010_00011_00000_100100	;
//memory[19]	<=	32'b000000_00001_00010_00011_00000_100100	;
//memory[20]	<=	32'b000000_00001_00010_00011_00000_100101	;
//memory[21]	<=	32'b000000_00001_00010_00011_00000_100101	;
//memory[22]	<=	32'b000000_00001_00010_00011_00000_100101	;
//memory[23]	<=	32'b000000_00001_00010_00011_00000_100101	;
//memory[24]	<=	32'b000000_00001_00010_00011_00000_100101	;
//memory[25]	<=	32'b000000_00001_00010_00011_00000_100101	;
//memory[26]	<=	32'b000000_00001_00010_00011_00000_100101	;
//memory[27]	<=	32'b000000_00001_00010_00011_00000_100101	;
//memory[28]	<=	32'b000000_00001_00010_00011_00000_100000	;
//memory[29]	<=	32'b000000_00001_00010_00011_00000_100000	;
//memory[30]	<=	32'b000000_00001_00010_00011_00000_100000	;
//memory[31]	<=	32'b000000_00001_00010_00011_00000_100000	;
//memory[32]	<=	32'b000000_00001_00010_00011_00000_100000	;
//memory[33]	<=	32'b000000_00001_00010_00011_00000_100000	;
//memory[34]	<=	32'b000000_00001_00010_00011_00000_100000	;
//memory[35]	<=	32'b000000_00001_00010_00011_00000_100000	;
//memory[36]	<=	32'b000000_00001_00010_00011_00000_100010	;
//memory[37]	<=	32'b000000_00001_00010_00011_00000_100010	;
//memory[38]	<=	32'b000000_00001_00010_00011_00000_100010	;
//memory[39]	<=	32'b000000_00001_00010_00011_00000_100010	;
//memory[40]	<=	32'b000000_00001_00010_00011_00000_100010	;
//memory[41]	<=	32'b000000_00001_00010_00011_00000_100010	;
//memory[42]	<=	32'b000000_00001_00010_00011_00000_100010	;
//memory[43]	<=	32'b000000_00001_00010_00011_00000_100010	;
//memory[44]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[45]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[46]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[47]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[48]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[49]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[50]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[51]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[52]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[53]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[54]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[55]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[56]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[57]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[58]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[59]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[60]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[61]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[62]	<=	32'b000000_00001_00001_00001_00000_100010	;
//memory[63]	<=	32'b000000_00001_00001_00001_00000_100010	;

//////// For IF
//
//memory[00]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[01]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[02]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[03]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[04]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[05]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[06]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[07]	<=	32'b000010_10101_10101_10101_10101_101010	;
//memory[08]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[09]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[10]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[11]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[12]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[13]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[14]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[15]	<=	32'b000000_00000_00000_00000_00000_000000	;
//

////// For MEM//////
//memory[00]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[01]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[02]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[03]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[04]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[05]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[06]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[07]	<=	32'b110011_10010_10011_10101_10101_101010	;
//memory[08]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[09]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[10]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[11]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[12]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[13]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[14]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[15]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[16]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[17]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[18]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[19]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[20]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[21]	<=	32'b000000_00000_00000_00000_00000_000000	;
//memory[22]	<=	32'b000000_00000_00000_00000_00000_000000	;



memory[00]	<=	32'b00000000000000000000000000000000	;
memory[01]	<=	32'b00000000000000000000000000000000	;
memory[02]	<=	32'b00000000000000000000000000000000	;
memory[03]	<=	32'b00000000000000000000000000000000	;
memory[04]	<=	32'b00000000000000000000000000000000	;
memory[05]	<=	32'b00000000000000000000000000000000	;
memory[06]	<=	32'b00000000000000000000000000000000	;
memory[07]	<=	32'b11001110010100111010110101101010	;
memory[08]	<=	32'b00000000000000000000000000000000	;
memory[09]	<=	32'b00000000000000000000000000000000	;
memory[10]	<=	32'b00000000000000000000000000000000	;
memory[11]	<=	32'b00000000000000000000000000000000	;
memory[12]	<=	32'b00000000000000000000000000000000	;
memory[13]	<=	32'b00000000000000000000000000000000	;
memory[14]	<=	32'b00000000000000000000000000000000	;
memory[15]	<=	32'b00000000000000000000000000000000	;

/////////////////////////////////////////////////////////
memory[16]	<=	32'b00000000001000010000100000100010	;
memory[17]	<=	32'b00000000000000000000000000000000	;
memory[18]	<=	32'b00000000000000000000000000000000	;
memory[19]	<=	32'b00000000000000000000000000000000	;
memory[20]	<=	32'b00000000000000000000000000000000	;
memory[21]	<=	32'b00000000000000000000000000000000	;
memory[22]	<=	32'b00000000000000000000000000000000	;
memory[23]	<=	32'b00010000001010011010000111110001	;
memory[24]	<=	32'b00000000000000000000000000000000	;
memory[25]	<=	32'b00000000000000000000000000000000	;
memory[26]	<=	32'b00000000000000000000000000000000	;
memory[27]	<=	32'b00000000000000000000000000000000	;
memory[28]	<=	32'b00000000000000000000000000000000	;
memory[29]	<=	32'b00000000000000000000000000000000	;
memory[30]	<=	32'b00000000000000000000000000000000	;
memory[31]	<=	32'b00000000000000000000000000000000	;


///////////////////////////////////////////////////////////
memory[32]	<=	32'b00111100001000011001101100110111	;
memory[33]	<=	32'b00111100010000100101011100101001	;
memory[34]	<=	32'b00000000000000000000000000000000	;
memory[35]	<=	32'b00000000000000000000000000000000	;
memory[36]	<=	32'b00000000000000000000000000000000	;
memory[37]	<=	32'b00000000000000000000000000000000	;
memory[38]	<=	32'b00000000000000000000000000000000	;
memory[39]	<=	32'b00000000000000000000000000000000	;
memory[40]	<=	32'b00000000000000000000000000000000	;
memory[41]	<=	32'b00000000001000100001100000100000	;
memory[42]	<=	32'b00000000001000100001100000100000	;
memory[43]	<=	32'b00000000001000100001100000100000	;
memory[44]	<=	32'b00000000001000100001100000100000	;
memory[45]	<=	32'b00000000001000100001100000100000	;
memory[46]	<=	32'b00000000001000100001100000100000	;
memory[47]	<=	32'b00000000000000000000000000000000	;
////////////////////////////////////////////////////////////////

memory[48]	<=	32'b00000000000000000000000000000000	;
memory[49]	<=	32'b00000000000000000000000000000000	;
memory[50]	<=	32'b00000000000000000000000000000000	;
memory[51]	<=	32'b00000000000000000000000000000000	;
memory[52]	<=	32'b00000000000000000000000000000000	;
memory[53]	<=	32'b00000000000000000000000000000000	;
memory[54]	<=	32'b00000000000000000000000000000000	;
memory[55]	<=	32'b10101100001100001010110101101010	;
memory[56]	<=	32'b10101100001100001010110101101010	;
memory[57]	<=	32'b10101100001100001010110101101010	;
memory[58]	<=	32'b10101100001100001010110101101010	;
memory[59]	<=	32'b10101100001100001010110101101010	;
memory[60]	<=	32'b10101100001100001010110101101010	;
memory[61]	<=	32'b00000000000000000000000000000000	;
memory[62]	<=	32'b00000000000000000000000000000000	;
memory[63]	<=	32'b00000000000000000000000000000000	;



	end
  
	dlx DLX(
	.PHI1	(clk),
	.DIn	(DIn),
	.IIn	(IIn),
	.MRST	(~MRST),
	.TCE	(`LogicZero),
	.TMS	(`LogicZero),
	.TDI	(`LogicZero),
	.DAddr	(DAddr),
	.DRead	(DRead),
	.DWrite	(DWrite),
	.DOut	(DOut),
	.IAddr	(IAddr),
	.IRead	(IRead),
	.TDO	(),
	.troout(troout)
	);

endmodule
